`include "icezum_adc.v"

module icezum_adc_tb;




endmodule
