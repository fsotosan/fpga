`include "ads7924.v"

module ads7924_tb;




endmodule
